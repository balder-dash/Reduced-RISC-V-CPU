module control #(
    parameters
) (
    input logic EQ,
    input logic instr, //needs unknown width
    output logic RegWrite,
    output logic ALUctrl,
    output logic ALUsrc,
    output logic ImmSrc,
    output logic PCsrc 
);
    
endmodule